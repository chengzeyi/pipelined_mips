`include "ctrl_encode_def.v"

module IF_ID_REG(clk, id_ex_flush, instruction_in);